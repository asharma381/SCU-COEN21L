module s1f0(a1, b1, F);
	input a1, b1;
	output F;
	
	assign F = a1^b1;
endmodule