module sum0(a0, b0, F);
	input a0, b0;
	output F;
	
	assign F = a0^b0;
endmodule